library IEEE;
use IEEE.std_logic_1164.all;

entity cpu is
	port (clock, reset : in std_logic;
		from_memory : in std_logic_vector (7 downto 0);
		write : out std_logic;
		address : out std_logic_vector (7 downto 0);
		to_memory : out std_logic_vector (7 downto 0));
end entity;

architecture cpu_arch of cpu is

	component control_unit
		port (clock, reset : in std_logic;
			IR : in std_logic_vector (7 downto 0);
			CCR_Result : in std_logic_vector (3 downto 0);
			IR_Load : out std_logic;
			MAR_Load : out std_logic;
			PC_Load : out std_logic;
			PC_Inc : out std_logic;
			A_Load : out std_logic;
			B_Load : out std_logic;
			ALU_Sel : out std_logic (2 downto 0);
			CCR_Load : out std_logic;
			Bus1_Sel : out std_logic_vector (1 downto 0);
			Bus2_Sel : out std_logic_vector (1 downto 0);
			write : out std_logic);
	end component;

	component data_path
		port (clock, reset : in std_logic;
			IR_Load : in std_logic;
			MAR_Load : in std_logic;
			PC_Load : in std_logic;
			PC_Inc : in std_logic;
			A_Load : in std_logic;
			B_Load : in std_logic;
			ALU_Sel : in std_logic_vector (2 downto 0);
			CCR_Load : in std_logic;
			Bus1_Sel : in std_logic_vector (1 downto 0);
			Bus2_Sel : in std_logic_vector (1 downto 0);
			from_memory : in std_logic_vector (7 downto 0);
			IR : out std_logic_vector (7 downto 0);
			CCR_Result : out std_logic_vector (3 downto 0);
			to_memory : out std_logic_vector (7 downto 0);
			address : out std_logic_vector (7 downto 0));
	end component;
			

	begin

end architecture;
